module ALU181(
  input [3:0] A,
  input [3:0] B,
  input C0,
  input M,  
  input [3:0] S,
  output reg C4,
  output reg [3:0] F,
  output AequB,
  output P,
  output G
  );
    always@(A or B or S or M or C0)
	begin
      case({S,M,C0})
        6'b0000_0_1: {C4, F} = A;
        6'b0000_0_0: {C4, F} = A+1;        
        6'b0000_1_1, 
        6'b0000_1_0: {C4, F} = {!A[3], !A[2], !A[1], !A[0]};       

        6'b0001_0_1: {C4, F} = A|B;
        6'b0001_0_0: {C4, F} = (A|B)+1;        
        6'b0001_1_1, 
        6'b0001_1_0: {C4, F} = ~(A|B);        

        6'b0010_0_1: {C4, F} = A|({!B[3], !B[2], !B[1], !B[0]});
        6'b0010_0_0: {C4, F} = (A|({!B[3], !B[2], !B[1], !B[0]}))+1;        
        6'b0010_1_1, 
        6'b0010_1_0: {C4, F} = ({!A[3], !A[2], !A[1], !A[0]})&B;        

        6'b0011_0_1: {C4, F} = 5'b01111;
        6'b0011_0_0: {C4, F} = 5'b10000;        
        6'b0011_1_1, 
        6'b0011_1_0: {C4, F} = 5'b00000;        

        6'b0100_0_1: {C4, F} = A+(A&({!B[3], !B[2], !B[1], !B[0]}));
        6'b0100_0_0: {C4, F} = (A+(A&({!B[3], !B[2], !B[1], !B[0]})))+1;        
        6'b0100_1_1, 
        6'b0100_1_0: {C4, F} = ~(A&B);        

        6'b0101_0_1: {C4, F} = (A&({!B[3], !B[2], !B[1], !B[0]}))+(A|B);
        6'b0101_0_0: {C4, F} = ((A&({!B[3], !B[2], !B[1], !B[0]}))+(A|B))+1;        
        6'b0101_1_1, 
        6'b0101_1_0: {C4, F} = {!B[3], !B[2], !B[1], !B[0]};        

        6'b0110_0_1: begin
						{C4, F} = A-B+5'b11111;
						C4=!C4;
					 end
        6'b0110_0_0: begin
						{C4, F} = A-B;
						C4=!C4; 
					 end
        6'b0110_1_1, 
        6'b0110_1_0: {C4, F} = A^B;        

        6'b0111_0_1: begin
						{C4, F} = (A&({!B[3], !B[2], !B[1], !B[0]}))+5'b11111;
						C4 = ~C4;
					 end
        6'b0111_0_0: begin
						{C4, F} = (A&({!B[3], !B[2], !B[1], !B[0]}));
						C4 = ~C4;
					 end
        6'b0111_1_1, 
        6'b0111_1_0: {C4, F} = (A&({!B[3], !B[2], !B[1], !B[0]}));        

        6'b1000_0_1: {C4, F} = A+(A&B);
        6'b1000_0_0: {C4, F} = A+(A&B)+1;        
        6'b1000_1_1, 
        6'b1000_1_0: {C4, F} = ({!A[3], !A[2], !A[1], !A[0]}|B);        

        6'b1001_0_1: {C4, F} = A+B;
        6'b1001_0_0: {C4, F} = A+B+1;        
        6'b1001_1_1, 
        6'b1001_1_0: {C4, F} = ~(A^B);        

        6'b1010_0_1: {C4, F} = (A&B)+(A|({!B[3], !B[2], !B[1], !B[0]}));
        6'b1010_0_0: {C4, F} = (A&B)+(A|({!B[3], !B[2], !B[1], !B[0]}))+1;        
        6'b1010_1_1, 
        6'b1010_1_0: {C4, F} = B;        

        6'b1011_0_1: begin
						{C4, F} = A&B+5'b11111;
						C4 = ~C4;
					 end
        6'b1011_0_0: begin
						{C4, F} = A&B; 
						C4 = ~C4;
					 end
        6'b1011_1_1, 
        6'b1011_1_0: {C4, F} = A&B;        

        6'b1100_0_1: {C4, F} = A+A;
        6'b1100_0_0: {C4, F} = A+A+1;        
        6'b1100_1_1, 
        6'b1100_1_0: {C4, F} = 4'b1111; //逻辑1       

        6'b1101_0_1: {C4, F} = A+(A|B);
        6'b1101_0_0: {C4, F} = A+(A|B)+1;        
        6'b1101_1_1, 
        6'b1101_1_0: {C4, F} = A|({!B[3], !B[2], !B[1], !B[0]});        

        6'b1110_0_1: {C4, F} = A+(A|({!B[3], !B[2], !B[1], !B[0]}));
        6'b1110_0_0: {C4, F} = A+(A|({!B[3], !B[2], !B[1], !B[0]}))+1;        
        6'b1110_1_1, 
        6'b1110_1_0: {C4, F} = A|B;        

        6'b1111_0_1: begin
						{C4, F} = A+5'b11111;
						C4 = ~C4;
					 end
        6'b1111_0_0: begin
						{C4, F} = A;
						C4 = ~C4;
					 end
        6'b1111_1_1, 
        6'b1111_1_0: {C4, F} = A;        
      endcase
	  C4 = ~C4;
	end
    assign AequB = F[0]&F[1]&F[2]&F[3];
	assign P=(A[0]^B[0])&(A[1]^B[1])&(A[2]^B[2])&(A[3]^B[3]);
	assign G=(A[3]&B[3])+(A[2]&B[2])&(A[3]^B[3])+(A[1]&B[1])&(A[2]^B[2])&(A[3]^B[3])+(A[0]&B[0])&(A[1]^B[1])&(A[2]^B[2])&(A[3]^B[3]); 
endmodule



